`include "opcodes.v"

module ID_EX(Clk, Reset_N);
    
endmodule